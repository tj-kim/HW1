// Simple Verilog test
module hello_test ();
initial begin
	$display("Hello, Comparch!");
end
endmodule